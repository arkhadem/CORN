library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE WORK.NewTypes.ALL;

ENTITY Neuron_Weights IS
    PORT(
        Clk : IN STD_LOGIC;
		Rst : IN STD_LOGIC;
        En : IN DecodedSelectorType;
        ADDR : IN  STD_LOGIC_VECTOR((LOGK - 1) DOWNTO 0);
        DATA : out InputWeightType
    );
END Neuron_Weights;

architecture Behavioral of Neuron_Weights is
    SIGNAL ROM: WeightMatrixType;
    SIGNAL rdata: InputWeightType;
begin
	process (Clk)
    begin
        if (Clk'event and Clk = '1') then
			if (Rst = '1') then
				ROM <= (
					("0000000000011100", "0000000001000010", "0000000000110011", "0000000001100000", "0000000001011101", "0000000001001010", "0000000010000111", "0000000001101101", "0000000010001000", "0000000001101001", "0000000011100001", "0000000001101101", "0000000001100000", "0000000010100011", "0000000001010010", "0000000011011000"),
					("0000000011000110", "0000000010101011", "0000000010001111", "0000000000001100", "0000000001101100", "0000000001001111", "0000000001000101", "0000000010001111", "0000000011110111", "0000000010000111", "0000000001001110", "0000000000110110", "0000000011001111", "0000000001101011", "0000000011100111", "0000000010000111"),
					("0000000001110111", "0000000001101110", "0000000010100110", "0000000000011001", "0000000011011000", "0000000011010100", "0000000001011111", "0000000001100000", "0000000010001011", "0000000011100101", "0000000010001010", "0000000000001110", "0000000010011000", "0000000010101110", "0000000000000111", "0000000010000000"),
					("0000000010010101", "0000000001101011", "0000000001111101", "0000000001001010", "0000000011100101", "0000000011100100", "0000000000001101", "0000000010110010", "0000000010010011", "0000000001011011", "0000000000000110", "0000000010000110", "0000000010110011", "0000000011011101", "0000000000001010", "0000000011001101"),
					("0000000000111100", "0000000010100001", "0000000001110100", "0000000010000011", "0000000001010010", "0000000011101010", "0000000010010001", "0000000010110110", "0000000001010000", "0000000010011110", "0000000011100110", "0000000010000111", "0000000010011110", "0000000011110110", "0000000011100011", "0000000011010011"),
					("0000000010000100", "0000000011100101", "0000000010001110", "0000000001000111", "0000000001011110", "0000000011011111", "0000000011100000", "0000000001000101", "0000000001010010", "0000000010110001", "0000000000000000", "0000000010000010", "0000000011000001", "0000000001000100", "0000000010110111", "0000000001010010"),
					("0000000000111110", "0000000001000000", "0000000011001110", "0000000011100100", "0000000011010011", "0000000000010001", "0000000011111100", "0000000011000100", "0000000000001010", "0000000001010011", "0000000001101101", "0000000001001000", "0000000000011100", "0000000011101000", "0000000000110010", "0000000011001110"),
					("0000000001010000", "0000000000101000", "0000000010101000", "0000000010001011", "0000000000011101", "0000000010010111", "0000000000110010", "0000000001010111", "0000000001011010", "0000000001001101", "0000000000110100", "0000000001000100", "0000000001111101", "0000000010100000", "0000000001011111", "0000000011101110")
				);
			end if;
		end if;
	end process;

    SINKS: for index in (N - 1) downto 0 generate
	begin
		SINK: rdata(index) <= ROM(index)(conv_integer(ADDR));
	end generate;

    process (Clk)
    begin
        if (Clk'event and Clk = '1') then
            for index in (N - 1) downto 0 loop
                if (En(index) = '1') then
                    DATA(index) <= rdata(index);
                end if;
            end loop;
        end if;
    end process;

end Behavioral;
